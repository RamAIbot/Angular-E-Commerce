package decode_test_pkg;
    import uvm_pkg::*;
    import uvmf_base_pkg::*; // IMPORTANT for uvmf_test_base
    import uvmf_base_pkg_hdl::*;
    import decode_env_pkg::*;
    import decode_in_pkg::*;
    import decode_out_pkg::*;

    `include "uvm_macros.svh"
    `include "src/print_component.svh"
    `include "src/test_top.svh"
    
    
endpackage